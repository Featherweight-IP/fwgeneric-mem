
/****************************************************************************
 * fwgeneric_sram_byte_en.v
 ****************************************************************************/

  
/**
 * Module: fwgeneric_sram_byte_en
 * 
 * TODO: Add module documentation
 */
module fwgeneric_sram_byte_en;


endmodule


